library verilog;
use verilog.vl_types.all;
entity Time_vlg_check_tst is
    port(
        t               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Time_vlg_check_tst;
