library verilog;
use verilog.vl_types.all;
entity Bcd_vlg_vec_tst is
end Bcd_vlg_vec_tst;
