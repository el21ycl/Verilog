library verilog;
use verilog.vl_types.all;
entity Bcd7seg_0_vlg_vec_tst is
end Bcd7seg_0_vlg_vec_tst;
