library verilog;
use verilog.vl_types.all;
entity Random_vlg_vec_tst is
end Random_vlg_vec_tst;
