library verilog;
use verilog.vl_types.all;
entity Key_vlg_vec_tst is
end Key_vlg_vec_tst;
